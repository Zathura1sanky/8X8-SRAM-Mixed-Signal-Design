* E:\FOSSEE\eSim\library\SubcircuitLibrary\Sanket_SRAM_CELL\Sanket_SRAM_CELL.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/04/22 13:31:57

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC3  Net-_SC1-Pad3_ Net-_SC2-Pad2_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC5  Net-_SC2-Pad2_ Net-_SC1-Pad3_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ GND sky130_fd_pr__nfet_01v8_lvt		
SC6  Net-_SC6-Pad1_ Net-_SC1-Pad2_ Net-_SC2-Pad2_ GND sky130_fd_pr__nfet_01v8_lvt		
SC2  Net-_SC1-Pad3_ Net-_SC2-Pad2_ Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
SC4  Net-_SC2-Pad2_ Net-_SC1-Pad3_ Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
U1  Net-_SC1-Pad1_ Net-_SC1-Pad3_ Net-_SC2-Pad3_ Net-_SC1-Pad2_ Net-_SC6-Pad1_ PORT		

.end
