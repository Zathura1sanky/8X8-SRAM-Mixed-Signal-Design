* E:\FOSSEE\ws\3x8DECODER_TEST\3x8DECODER_TEST.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/05/22 17:32:35

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  a2 a1 a0 Net-_U5-Pad4_ Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_4		
U6  Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad8_ Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ y7 y6 y5 y4 y3 y2 y1 y0 dac_bridge_8		
v4  Net-_U5-Pad4_ GND DC		
v3  a0 GND pulse		
v2  a1 GND pulse		
v1  a2 GND pulse		
U9  y5 plot_v1		
U10  y4 plot_v1		
U7  y7 plot_v1		
U8  y6 plot_v1		
U11  y3 plot_v1		
U12  y2 plot_v1		
U13  y1 plot_v1		
U14  y0 plot_v1		
U1  a2 plot_v1		
U2  a1 plot_v1		
U4  a0 plot_v1		
scmode1  SKY130mode		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad8_ Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ sanket_decoder_3x8		

.end
