* E:\FOSSEE\eSim\library\SubcircuitLibrary\BIT_ADDRESSABLE_SRAM_1BIT\BIT_ADDRESSABLE_SRAM_1BIT.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/07/22 17:52:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U4-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ SANKET_1BIT_SRAM		
U3  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U4  Net-_U1-Pad3_ Net-_U4-Pad2_ dac_bridge_1		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ PORT		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ ? sanket_write_ckt		

.end
